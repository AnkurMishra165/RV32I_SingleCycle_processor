// data_mem.v - data memory
module data_mem #(parameter DATA_WIDTH = 32, ADDR_WIDTH = 32, MEM_SIZE = 64) (
    input                     clk,
    input                     wr_en,
    input       [2:0]         funct3,
    input       [ADDR_WIDTH-1:0] wr_addr,
    input       [DATA_WIDTH-1:0] wr_data,
    output reg  [DATA_WIDTH-1:0] rd_data_mem
);

  // 64 x 32-bit words
  reg [DATA_WIDTH-1:0] data_ram [0:MEM_SIZE-1];

  // word index (use ADDR_WIDTH for slicing; addresses are byte-addressed)
  wire [ADDR_WIDTH-1:0] word_addr = wr_addr[ADDR_WIDTH-1:2] % MEM_SIZE;

  // =======================
  // Synchronous WRITE path
  // =======================
  always @(posedge clk) begin
    if (wr_en) begin
      case (funct3)
        3'b000: begin // SB
          case (wr_addr[1:0])
            2'b00: data_ram[word_addr][7:0]   <= wr_data[7:0];
            2'b01: data_ram[word_addr][15:8]  <= wr_data[7:0];
            2'b10: data_ram[word_addr][23:16] <= wr_data[7:0];
            2'b11: data_ram[word_addr][31:24] <= wr_data[7:0];
          endcase
        end

        3'b001: begin // SH  
          if (wr_addr[1] == 1'b0) begin
            // lower halfword (bits [15:0])
            data_ram[word_addr][15:0] <= wr_data[15:0];
          end else begin
            // upper halfword (bits [31:16])
            data_ram[word_addr][31:16] <= wr_data[15:0];
          end
        end

        3'b010: begin // SW
          data_ram[word_addr] <= wr_data;
        end
        default: ; // no store
      endcase
    end
  end

  // ======================
  // Combinational READ path
  // ======================
  always @(*) begin
    case (funct3)
      3'b000: begin // LB
        case (wr_addr[1:0])
          2'b00: rd_data_mem = {{24{data_ram[word_addr][7]}},   data_ram[word_addr][7:0]};
          2'b01: rd_data_mem = {{24{data_ram[word_addr][15]}},  data_ram[word_addr][15:8]};
          2'b10: rd_data_mem = {{24{data_ram[word_addr][23]}},  data_ram[word_addr][23:16]};
          2'b11: rd_data_mem = {{24{data_ram[word_addr][31]}},  data_ram[word_addr][31:24]};
        endcase
      end

      3'b001: begin // LH  
        if (wr_addr[1] == 1'b0) begin
          rd_data_mem = {{16{data_ram[word_addr][15]}}, data_ram[word_addr][15:0]};
        end else begin
          rd_data_mem = {{16{data_ram[word_addr][31]}}, data_ram[word_addr][31:16]};
        end
      end

      3'b010: begin // LW
        rd_data_mem = data_ram[word_addr];
      end

      3'b100: begin // LBU
        case (wr_addr[1:0])
          2'b00: rd_data_mem = {24'b0, data_ram[word_addr][7:0]};
          2'b01: rd_data_mem = {24'b0, data_ram[word_addr][15:8]};
          2'b10: rd_data_mem = {24'b0, data_ram[word_addr][23:16]};
          2'b11: rd_data_mem = {24'b0, data_ram[word_addr][31:24]};
        endcase
      end

      3'b101: begin // LHU  
        if (wr_addr[1] == 1'b0)
          rd_data_mem = {16'b0, data_ram[word_addr][15:0]};
        else
          rd_data_mem = {16'b0, data_ram[word_addr][31:16]};
      end

      default: rd_data_mem = 32'b0;
    endcase
  end

endmodule


